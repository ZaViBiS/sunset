module config

pub const url = 'https://api.sunrise-sunset.org/json?lat=48.501792&lng=35.060611&formatted=0&date='
pub const today_url = url + 'today'
pub const tomorrow_url = url + 'tomorrow'
pub const blynk_url = 'http://blynk.cloud/external/api/batch/update?token=sq-8rXjk0R4pfAqxjF1XCNaxbMFHkPm_&d0='
pub const error_time = '2021-01-01 00:00:00'
pub const art = '                          _   
 ___ _   _ _ __  ___  ___| |_ 
/ __| | | | \'_ \\/ __|/ _ \\ __|
\\__ \\ |_| | | | \\__ \\  __/ |_ 
|___/\\__,_|_| |_|___/\\___|\\__|
                            '
